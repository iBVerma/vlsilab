module xor_gate (
    input clk,
    input a,
    input b,
    output y
);

assign y = a ^ b;

endmodule
